module obj

pub enum LogLevel {
	debug = 0
	information = 1
	log = 2
	warn = 3
	error = 4
	fatal = 5
}
