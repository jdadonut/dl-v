module obj

pub enum Services {
	gelbooru
	danbooru
	safebooru
}
