module obj

enum services {
	Gelbooru
	Danbooru
	Safebooru
}