module util
// fn XML.parseAttrsFromNodeType() {
// 	// <string .*?name="file_url".*?>(.+)</string>
// }
// fn XML.parseNodes() {
// 	// <primaryAddress.*>((.|\n)*?)<\/primaryAddress>
// }