module obj

enum logLevel {
	DEBUG
	INFORMATION
	LOG
	WARN
	ERROR
	FATAL
}
